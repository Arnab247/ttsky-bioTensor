`default_nettype none

module norm_seed_lut (
    input  wire [31:0] d_in,    // Always 1.0 to 1.999 (Q16.16)
    output reg  [31:0] seed_out // Guesses 0.5 to 1.0 (Q16.16)
);
    // Look at the top 5 bits of the fraction (bits 15:11)
    wire [4:0] index = d_in[15:11];

    always @(*) begin
        case (index)
            // Pre-calculated 1/x for the range [1.0, 2.0)
            5'd0:  seed_out = 32'h0000_FE00; // 1 / 1.015 = 0.985
            5'd1:  seed_out = 32'h0000_F400; // 1 / 1.046 = 0.953
            5'd2:  seed_out = 32'h0000_EB00; // 1 / 1.078 = 0.917
            5'd3:  seed_out = 32'h0000_E200; // 1 / 1.109 = 0.882
            5'd4:  seed_out = 32'h0000_DA00; // 1 / 1.140 = 0.851
            5'd5:  seed_out = 32'h0000_D200; // 1 / 1.171 = 0.820
            5'd6:  seed_out = 32'h0000_CB00; // 1 / 1.203 = 0.792
            5'd7:  seed_out = 32'h0000_C400; // 1 / 1.234 = 0.765
            5'd8:  seed_out = 32'h0000_BE00; // 1 / 1.265 = 0.742
            5'd9:  seed_out = 32'h0000_B800; // 1 / 1.296 = 0.718
            5'd10: seed_out = 32'h0000_B200; // 1 / 1.328 = 0.695
            5'd11: seed_out = 32'h0000_AC00; // 1 / 1.359 = 0.671
            5'd12: seed_out = 32'h0000_A700; // 1 / 1.390 = 0.652
            5'd13: seed_out = 32'h0000_A200; // 1 / 1.421 = 0.632
            5'd14: seed_out = 32'h0000_9E00; // 1 / 1.453 = 0.617
            5'd15: seed_out = 32'h0000_9900; // 1 / 1.484 = 0.597
            5'd16: seed_out = 32'h0000_9500; // 1 / 1.515 = 0.582
            5'd17: seed_out = 32'h0000_9100; // 1 / 1.546 = 0.566
            5'd18: seed_out = 32'h0000_8D00; // 1 / 1.578 = 0.550
            5'd19: seed_out = 32'h0000_8900; // 1 / 1.609 = 0.535
            5'd20: seed_out = 32'h0000_8600; // 1 / 1.640 = 0.523
            5'd21: seed_out = 32'h0000_8300; // 1 / 1.671 = 0.511
            5'd22: seed_out = 32'h0000_8000; // 1 / 1.703 = 0.500
            5'd23: seed_out = 32'h0000_7D00; // 1 / 1.734 = 0.488
            5'd24: seed_out = 32'h0000_7A00; // 1 / 1.765 = 0.476
            5'd25: seed_out = 32'h0000_7800; // 1 / 1.796 = 0.468
            5'd26: seed_out = 32'h0000_7500; // 1 / 1.828 = 0.457
            5'd27: seed_out = 32'h0000_7300; // 1 / 1.859 = 0.449
            5'd28: seed_out = 32'h0000_7100; // 1 / 1.890 = 0.441
            5'd29: seed_out = 32'h0000_6E00; // 1 / 1.921 = 0.429
            5'd30: seed_out = 32'h0000_6C00; // 1 / 1.953 = 0.421
            5'd31: seed_out = 32'h0000_6A00; // 1 / 1.984 = 0.414
        endcase
    end
endmodule